library ieee;
USE ieee.std_logic_1164.all;

ENTITY Exp4b IS
  PORT (SW: IN STD_LOGIC_VECTOR(17 downto 0);
		HEX0: OUT STD_LOGIC_VECTOR(0 to 6);
		HEX1: OUT STD_LOGIC_VECTOR(0 to 6);		
		HEX2: OUT STD_LOGIC_VECTOR(0 to 6);
		HEX3: OUT STD_LOGIC_VECTOR(0 to 6);
		--HEX4: OUT STD_LOGIC_VECTOR(0 to 6);
		--HEX5: OUT STD_LOGIC_VECTOR(0 to 6);
		--HEX6: OUT STD_LOGIC_VECTOR(0 to 6);
		--HEX7: OUT STD_LOGIC_VECTOR(0 to 6);
		LEDR: OUT STD_LOGIC_VECTOR(17 downto 0);
		KEY : IN STD_LOGIC_VECTOR(3 downto 0));
END Exp4b;

ARCHITECTURE experimento OF Exp4b IS
	
	COMPONENT Contador IS
	  PORT (enb, clk, clr : IN STD_LOGIC ;
		  Q : OUT STD_LOGIC_VECTOR(15 downto 0));
	END COMPONENT Contador;
	
	COMPONENT Decoder IS
		PORT (s: in std_logic_vector(3 downto 0);
			b: out std_logic_vector(0 to 6));
	END COMPONENT Decoder;
	
	SIGNAL Nclock : STD_LOGIC;
	SIGNAL Nclear : STD_LOGIC;
	SIGNAL Q : STD_LOGIC_VECTOR(15 downto 0);
	SIGNAL Nenable : STD_LOGIC;
	
	BEGIN
	Nclock <= NOT KEY(0);
	Nclear <= NOT KEY(1);
	
	
	B01 : Contador port map(KEY(2), Nclock, Nclear, Q);
	B02 : Decoder port map (Q(3 downto 0), HEX0(0 to 6));
	B03 : Decoder port map (Q(7 downto 4), HEX1(0 to 6));
	B04 : Decoder port map (Q(11 downto 8), HEX2(0 to 6));
	B05 : Decoder port map (Q(15 downto 12), HEX3(0 to 6));
	
	LEDR(15 downto 0) <= Q;
	
	
END experimento;